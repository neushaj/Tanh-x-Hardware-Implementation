library verilog;
use verilog.vl_types.all;
entity PartD_Q_TB is
end PartD_Q_TB;
