library verilog;
use verilog.vl_types.all;
entity PartD_TB is
end PartD_TB;
