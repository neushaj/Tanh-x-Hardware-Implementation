library verilog;
use verilog.vl_types.all;
entity adder is
    port(
        A               : in     vl_logic_vector(15 downto 0);
        B               : in     vl_logic_vector(15 downto 0);
        sub_sel         : in     vl_logic;
        R               : out    vl_logic_vector(15 downto 0)
    );
end adder;
