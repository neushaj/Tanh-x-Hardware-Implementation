library verilog;
use verilog.vl_types.all;
entity PartF_TB is
end PartF_TB;
